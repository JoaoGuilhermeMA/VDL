library verilog;
use verilog.vl_types.all;
entity grayJohnson_vlg_vec_tst is
end grayJohnson_vlg_vec_tst;
