library verilog;
use verilog.vl_types.all;
entity paridadePar_vlg_vec_tst is
end paridadePar_vlg_vec_tst;
