library verilog;
use verilog.vl_types.all;
entity paridadePar_vlg_check_tst is
    port(
        saida           : in     vl_logic_vector(0 to 1);
        sampler_rx      : in     vl_logic
    );
end paridadePar_vlg_check_tst;
