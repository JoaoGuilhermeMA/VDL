library verilog;
use verilog.vl_types.all;
entity acionamentoMaquinas_vlg_vec_tst is
end acionamentoMaquinas_vlg_vec_tst;
