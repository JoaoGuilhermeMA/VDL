library verilog;
use verilog.vl_types.all;
entity acionamentoMaquinas_vlg_check_tst is
    port(
        m1              : in     vl_logic;
        m2              : in     vl_logic;
        m3              : in     vl_logic;
        m4              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end acionamentoMaquinas_vlg_check_tst;
