library verilog;
use verilog.vl_types.all;
entity BCDDoisEntreCinco_vlg_vec_tst is
end BCDDoisEntreCinco_vlg_vec_tst;
